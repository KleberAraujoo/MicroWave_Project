`timescale 1s/1ns
`include "controler.v"

module controler_tb();

    reg startn, stopn, clearn, door_closed, clock;
    reg [9:0] keypad;
    wire mag_on;
    wire[6:0] sec_ones_segs, sec_tens_segs, mins_segs;

    controler DUT(
        .startn(startn),
        .stopn(stopn),
        .clearn(clearn),
        .door_closed(door_closed),
        .clock(clock),
        .keypad(keypad),
        .mag_on(mag_on),
        .sec_ones_segs(sec_ones_segs),
        .sec_tens_segs(sec_tens_segs),
        .mins_segs(mins_segs)
        );

    initial clock = 0;

    //parameter secs = 1000;
    parameter Wait = 0.5;

    always #0.005 clock = ~clock;

    initial begin
        $dumpfile("controler_tb.vcd");
        $dumpvars(0, controler_tb);
    end

    initial begin

        keypad = 0; startn = 1; stopn = 1; clearn =1; door_closed = 1;

        //Caso 0: Funcionamento normal

        //Wait = 0.5;
        #(Wait) keypad = 1<< 1;
        #(Wait) keypad = 0;
        #(Wait) keypad = 1<< 3;
        #(Wait) keypad = 0;
        #(Wait) keypad = 1<< 0;
        #(Wait) keypad = 0;

        //Alguns casos podem ser testados durante o caso 0:

            //Caso 1: Tentar ligar com a porta aberta

            #(Wait) door_closed = 0;

            #(Wait) startn = 0;
            #(Wait) startn = 1;

            #(Wait) door_closed = 1;

            #(Wait) startn = 0;
            #(Wait) startn = 1;

            //Caso 2: Apertar start com microondas ligado

            #5 startn = 0;
            #(Wait) startn = 1;

            //Caso 3: abrir a porta com o microondas ligado

            #5 door_closed = 0;
            #5 door_closed = 1;

            #5 startn = 0;
            #(Wait) startn = 1;

            //Caso 4: apertar stop

            #5 stopn = 0;
            #5 stopn = 1;

            #5 startn = 0;
            #(Wait) startn = 1;


        #80;

        //Caso 5: Teste do Clear e tentar apertar dois botões quase que simultaneamente
        
        //Wait = 0.06;
        #(Wait);
        
        #(Wait) keypad = 1<< 8;
        #(Wait) keypad = 0;
        #(Wait) keypad = 1<< 5;
        #(Wait) keypad = 0;
        #(Wait) keypad = 1<< 1;
        #(Wait) keypad = 0;

        #(Wait) clearn = 0;
        #(Wait) clearn = 1;

        //5.1 Intervalo MAIOR que 4 bordas de relógio (40ms)

        #(Wait) keypad = 1<< 8;
        #(Wait) keypad = 0;
        #(Wait) keypad = 1<< 5;
        #(Wait) keypad = 10'b0000100010;
        #(Wait) keypad = 0;
        #(Wait);

        #(Wait) clearn = 0;
        #(Wait) clearn = 1;

        //5.2 Intervalo MENOR que 4 bordas de relógio (40ms)

        #(Wait) keypad = 1<< 8;
        #(Wait) keypad = 0;
        #(Wait) keypad = 1<< 5;
        #0.03   keypad = 10'b0000100010;
        #(Wait -0.03) keypad = 0;
        #(Wait);

        #(Wait) clearn = 0;
        #(Wait) clearn = 1;

        $finish();
    end




endmodule
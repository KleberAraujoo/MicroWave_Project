module seg7_driver (input wire [3:0] sec_ones, sec_tens, mins,
                                    output wire [6:0] sec_ones_segs, sec_tens_segs, mins_segs);


    assign sec_ones_segs = 
    /* 0 */ (sec_ones == 4'b0000) ? 7'b000_0001 : 
    /* 1 */ (sec_ones == 4'b0001) ? 7'b100_1111 :
    /* 2 */ (sec_ones == 4'b0010) ? 7'b001_0010 :
    /* 3 */ (sec_ones == 4'b0011) ? 7'b000_0110 :
    /* 4 */ (sec_ones == 4'b0100) ? 7'b100_1100 :
    /* 5 */ (sec_ones == 4'b0101) ? 7'b010_0100 :
    /* 6 */ (sec_ones == 4'b0110) ? 7'b010_0000 :
    /* 7 */ (sec_ones == 4'b0111) ? 7'b000_1111 :
    /* 8 */ (sec_ones == 4'b1000) ? 7'b000_0000 :
    /* 9 */ (sec_ones == 4'b1001) ? 7'b000_0100 :
    /* d */ 7'b000_0001;

        assign sec_tens_segs = 
    /* 0 */ (sec_tens == 4'b0000) ? 7'b000_0001 : 
    /* 1 */ (sec_tens == 4'b0001) ? 7'b100_1111 :
    /* 2 */ (sec_tens == 4'b0010) ? 7'b001_0010 :
    /* 3 */ (sec_tens == 4'b0011) ? 7'b000_0110 :
    /* 4 */ (sec_tens == 4'b0100) ? 7'b100_1100 :
    /* 5 */ (sec_tens == 4'b0101) ? 7'b010_0100 :
    /* 6 */ (sec_tens == 4'b0110) ? 7'b010_0000 :
    /* 7 */ (sec_tens == 4'b0111) ? 7'b000_1111 :
    /* 8 */ (sec_tens == 4'b1000) ? 7'b000_0000 :
    /* 9 */ (sec_tens == 4'b1001) ? 7'b000_0100 :
    /* d */ 7'b000_0001;

    assign mins_segs = 
    /* 0 */ (mins == 4'b0000) ? 7'b000_0001 : 
    /* 1 */ (mins == 4'b0001) ? 7'b100_1111 :
    /* 2 */ (mins == 4'b0010) ? 7'b001_0010 :
    /* 3 */ (mins == 4'b0011) ? 7'b000_0110 :
    /* 4 */ (mins == 4'b0100) ? 7'b100_1100 :
    /* 5 */ (mins == 4'b0101) ? 7'b010_0100 :
    /* 6 */ (mins == 4'b0110) ? 7'b010_0000 :
    /* 7 */ (mins == 4'b0111) ? 7'b000_1111 :
    /* 8 */ (mins == 4'b1000) ? 7'b000_0000 :
    /* 9 */ (mins == 4'b1001) ? 7'b000_0100 :
    /* d */ 7'b000_0001;

    
endmodule